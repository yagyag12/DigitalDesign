`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.03.2024 12:45:55
// Design Name: 
// Module Name: Display7seg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Display7seg(
    input wire [3:0] A,
    output wire [6:0] Y,
    output wire DP,
    output wire [7:0] AN
    );
    
    assign AN = 8'b11111110;
    assign DP = 1'b1;
    
    assign Y[0] = (~A[3] && ~A[2] && ~A[1] && A[0]) | (~A[3] && A[2] && ~A[1] && ~A[0]) 
                    | (A[3] && ~A[2] && A[1] && A[0]) | (A[3] && A[2] && ~A[1] && A[0]);
                    
    assign Y[1] = (~A[3] && A[2] && ~A[1] && A[0]) | (~A[3] && A[2] && A[1] && ~A[0]) |
                    (A[3] && ~A[2] && A[1] && A[0]) | (A[3] && A[2] && ~A[1] && ~A[0]) |
                    (A[3] && A[2] && A[1] && ~A[0]) | (A[3] && A[2] && A[1] && A[0]);
                    
    assign Y[2] = (~A[3] && ~A[2] && A[1] && ~A[0]) | (A[3] && A[2] && ~A[1] && ~A[0]) |
                    (A[3] && A[2] && A[1] && ~A[0]) | (A[3] && A[2] && A[1] && A[0]);
                    
    assign Y[3] = (~A[3] && ~A[2] && ~A[1] && A[0]) | (~A[3] && A[2] && ~A[1] && ~A[0]) |
                    (~A[3] && A[2] && A[1] && A[0]) | (A[3] && ~A[2] && A[1] && ~A[0]) |
                    (A[3] && A[2] && A[1] && A[0]);
    
    assign Y[4] = (~A[3] && ~A[2] && ~A[1] && A[0]) | (~A[3] && ~A[2] && A[1] && A[0]) |
                    (~A[3] && A[2] && ~A[1] && ~A[0]) | (~A[3] && A[2] && ~A[1] && A[0]) |
                    (~A[3] && A[2] && A[1] && A[0]) | (A[3] && ~A[2] && ~A[1] && A[0]);
    
    assign Y[5] = (~A[3] && ~A[2] && ~A[1] && A[0]) | (~A[3] && ~A[2] && A[1] && ~A[0]) |
                    (~A[3] && ~A[2] && A[1] && A[0]) | (A[3] && A[2] && ~A[1] && A[0]);
                    
    assign Y[6] = (~A[3] && ~A[2] && ~A[1] && ~A[0]) | (~A[3] && ~A[2] && ~A[1] && A[0])|
                    (~A[3] && A[2] && A[1] && A[0]) | (A[3] && A[2] && ~A[1] && ~A[0]);

endmodule
